typedef struct {
    byte val1;
    int val2;
    string val3;
} data;